LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY multiplicador IS
PORT (
	A3 : IN std_logic;
	A2 : IN std_logic;
	A1 : IN std_logic;
	A0 : IN std_logic;
	B3 : IN std_logic;
	B2 : IN std_logic;
	B1 : IN std_logic;
	B0 : IN std_logic;
	S7 : OUT std_logic;
	S6 : OUT std_logic;
	S5 : OUT std_logic;
	S4 : OUT std_logic;
	S3 : OUT std_logic;
	S2 : OUT std_logic;
	S1 : OUT std_logic;
	S0 : OUT std_logic);
END multiplicador;

ARCHITECTURE data_flow OF multiplicador IS
BEGIN

S7 <= (A3 AND A1 AND A0 AND B3 AND B2) OR (A3 AND A2 AND A0 AND B3 AND B1) OR (A3 AND A1 AND B3 AND B2 AND B0) OR (A3 AND A2 AND B3
     AND B1 AND B0) OR (A3 AND A2 AND B3 AND B2) OR (A3 AND A2 AND A1 AND B3 AND B1) OR (A3 AND A1 AND B3 AND B2 AND B1) OR (A3
     AND A2 AND A1 AND A0 AND B3 AND B0) OR (A3 AND A0 AND B3 AND B2 AND B1 AND B0);

S6 <= (A2 AND A1 AND A0 AND B3 AND B2 AND B0) OR (A2 AND A0 AND B3 AND B2 AND B1 AND B0) OR (A2 AND A1 AND B3 AND B2 AND B1) OR (NOT A3
     AND A2 AND A1 AND B3 AND B2) OR (NOT A3 AND A2 AND A1 AND A0 AND B3 AND B1) OR (A3 AND A2 AND NOT B3 AND B2 AND B1) OR (A3 AND A1 AND A0
     AND NOT B3 AND B2 AND B1) OR (A3 AND A2 AND A0 AND NOT B3 AND B2 AND B0) OR (NOT A3 AND A2 AND A0 AND B3 AND B2 AND B0) OR (NOT A3 AND A2
     AND A1 AND B3 AND B1 AND B0) OR (A3 AND A1 AND NOT B3 AND B2 AND B1 AND B0) OR (NOT A3 AND A2 AND A0 AND B3 AND B2 AND B1) OR (A3 AND A2
     AND A1 AND NOT B3 AND B2 AND B0) OR (A3 AND NOT A2 AND B3 AND NOT B2) OR (A3 AND NOT A1 AND B3 AND NOT B2 AND NOT B1) OR (A3 AND NOT A2 AND NOT A1
     AND B3 AND NOT B1) OR (A3 AND B3 AND NOT B2 AND NOT B1 AND NOT B0) OR (A3 AND NOT A2 AND NOT A0 AND B3 AND NOT B1 AND NOT B0) OR (A3 AND NOT A1 AND NOT A0
     AND B3 AND NOT B2 AND NOT B0) OR (A3 AND NOT A2 AND NOT A1 AND B3 AND NOT B0) OR (A3 AND NOT A0 AND B3 AND NOT B2 AND NOT B1) OR (A3 AND NOT A2 AND NOT A1
     AND NOT A0 AND B3);

S5 <= (A3 AND A1 AND NOT A0 AND B2 AND NOT B1 AND NOT B0) OR (A2 AND NOT A1 AND NOT A0 AND B3 AND B1 AND NOT B0) OR (A2 AND NOT A0 AND B3 AND NOT B2 AND NOT B1) OR (
    NOT A3 AND A1 AND A0 AND B3 AND B2 AND B1) OR (A2 AND A1 AND NOT B3 AND B2 AND B1 AND B0) OR (A3 AND A2 AND A1 AND B2 AND NOT B1 AND NOT B0) OR (
    A3 AND A1 AND A0 AND B3 AND B1 AND B0) OR (A3 AND NOT A1 AND NOT A0 AND B3 AND B2 AND B1) OR (A3 AND A2 AND NOT A1 AND A0 AND B3 AND NOT B1 AND B0) OR (
    A3 AND NOT A2 AND NOT A1 AND B2 AND NOT B1) OR (A2 AND B3 AND NOT B2 AND NOT B1 AND NOT B0) OR (A3 AND A1 AND A0 AND NOT B2 AND B1 AND B0) OR (
    NOT A2 AND A1 AND A0 AND B3 AND B1 AND B0) OR (NOT A3 AND A2 AND A1 AND NOT B3 AND B2 AND B1) OR (NOT A3 AND A2 AND NOT A1 AND B3 AND NOT B2) OR (
    A3 AND NOT A2 AND NOT B3 AND B2 AND NOT B1) OR (NOT A3 AND A2 AND NOT A0 AND B3 AND NOT B2 AND NOT B0) OR (A3 AND NOT A2 AND NOT A0 AND NOT B3 AND B2 AND NOT B0) OR (
    NOT A3 AND A2 AND A1 AND A0 AND NOT B3 AND B2 AND B0) OR (NOT A3 AND A2 AND A0 AND NOT B3 AND B2 AND B1 AND B0) OR (NOT A3 AND NOT A2 AND A1 AND A0
     AND B3 AND B2) OR (A3 AND A2 AND NOT B3 AND NOT B2 AND B1 AND B0) OR (A3 AND NOT A2 AND A1 AND B3 AND NOT B2 AND B1) OR (NOT A3 AND A2 AND B3
     AND NOT B2 AND NOT B1) OR (A3 AND NOT A2 AND NOT A1 AND NOT B3 AND B2) OR (A3 AND NOT A2 AND A1 AND A0 AND B3 AND NOT B2 AND B0) OR (A3 AND NOT A2
     AND A0 AND B3 AND NOT B2 AND B1 AND B0) OR (A3 AND NOT B3 AND B2 AND NOT B1 AND NOT B0) OR (NOT A3 AND A2 AND NOT A1 AND NOT A0 AND B3) OR (NOT A3
     AND A2 AND NOT A1 AND B3 AND NOT B1 AND NOT B0) OR (A3 AND NOT A1 AND NOT A0 AND NOT B3 AND B2 AND NOT B1) OR (A3 AND NOT A1 AND B3 AND B2 AND B1 AND NOT B0) OR (
    A3 AND A2 AND A1 AND NOT A0 AND B3 AND NOT B1);

S4 <= (NOT A3 AND A1 AND A0 AND NOT B3 AND B2 AND B1 AND B0) OR (A2 AND NOT B3 AND B2 AND NOT B1 AND NOT B0) OR (NOT A3 AND A2 AND NOT A1 AND NOT A0 AND B2) OR (
    A3 AND A1 AND NOT A0 AND NOT B3 AND B1 AND NOT B0) OR (NOT A3 AND A1 AND NOT A0 AND B3 AND B1 AND NOT B0) OR (A3 AND A2 AND A1 AND A0 AND B1 AND NOT B0) OR (
    A1 AND NOT A0 AND B3 AND B2 AND B1 AND B0) OR (A2 AND NOT A1 AND B2 AND NOT B1 AND NOT B0) OR (A2 AND A0 AND B2 AND NOT B1 AND NOT B0) OR (A2
     AND NOT A1 AND NOT A0 AND B2 AND B0) OR (NOT A3 AND A1 AND B3 AND NOT B2 AND NOT B1) OR (A3 AND NOT A2 AND NOT A1 AND NOT B3 AND B1) OR (A3 AND NOT A1
     AND A0 AND B3 AND NOT B2 AND NOT B1 AND B0) OR (NOT A3 AND A2 AND NOT A1 AND NOT B3 AND B2 AND NOT B1) OR (NOT A3 AND A2 AND A1 AND NOT B3 AND NOT B2 AND B1
     AND B0) OR (NOT A3 AND NOT A2 AND A1 AND A0 AND NOT B3 AND B2 AND B1) OR (A3 AND NOT A2 AND A1 AND NOT B3 AND B2 AND NOT B1 AND B0) OR (NOT A3
     AND A2 AND NOT A1 AND A0 AND B3 AND NOT B2 AND B1) OR (A3 AND NOT A2 AND NOT A1 AND A0 AND B3 AND NOT B1 AND B0) OR (A3 AND NOT B3 AND NOT B2 AND B1 AND NOT B0) OR (
    NOT A3 AND NOT A2 AND A1 AND B3 AND NOT B2 AND NOT B0) OR (A3 AND NOT A2 AND NOT A0 AND NOT B3 AND NOT B2 AND B1) OR (NOT A3 AND NOT A2 AND A1 AND NOT A0 AND B3) OR (
    A1 AND B3 AND NOT B2 AND NOT B1 AND NOT B0) OR (A3 AND NOT A2 AND NOT A1 AND B1 AND NOT B0) OR (NOT A3 AND A2 AND NOT A1 AND NOT B3 AND B2 AND NOT B0) OR (
    A1 AND NOT A0 AND B3 AND NOT B2 AND NOT B1) OR (NOT A3 AND A2 AND NOT A0 AND NOT B3 AND B2 AND NOT B1) OR (A3 AND NOT A2 AND NOT A1 AND NOT A0 AND B1) OR (
    A3 AND NOT A2 AND A1 AND A0 AND B3 AND NOT B2 AND B1 AND B0) OR (NOT A3 AND A2 AND A1 AND A0 AND B3 AND NOT B1) OR (A3 AND NOT A1 AND NOT B3 AND B2
     AND B1 AND B0) OR (NOT A2 AND A1 AND NOT A0 AND B3 AND NOT B1 AND NOT B0) OR (A3 AND NOT A1 AND NOT A0 AND NOT B2 AND B1 AND NOT B0) OR (A3 AND A0
     AND B3 AND B2 AND B1 AND NOT B0) OR (A3 AND A2 AND A1 AND NOT A0 AND B3 AND B0);

S3 <= (A3 AND A2 AND NOT A1 AND B3 AND B2 AND NOT B1 AND B0) OR (A3 AND NOT A2 AND A1 AND B3 AND NOT B2 AND B1 AND B0) OR (A2 AND A0 AND NOT B3 AND B1
     AND NOT B0) OR (NOT A3 AND A0 AND B3 AND B2 AND B1 AND B0) OR (NOT A3 AND A1 AND NOT A0 AND B2 AND B0) OR (A3 AND A2 AND A1 AND A0 AND NOT B3
     AND B0) OR (NOT A2 AND A0 AND B3 AND B1 AND NOT B0) OR (A3 AND A1 AND NOT A0 AND NOT B2 AND B0) OR (A0 AND B3 AND NOT B2 AND NOT B1 AND NOT B0) OR (
    A1 AND NOT A0 AND B2 AND NOT B1 AND NOT B0) OR (A1 AND NOT B3 AND B2 AND NOT B1 AND NOT B0) OR (NOT A3 AND NOT A2 AND NOT A1 AND A0 AND B3) OR (NOT A3
     AND A2 AND NOT A1 AND NOT A0 AND B1) OR (A3 AND NOT A2 AND NOT A1 AND NOT B3 AND B0) OR (NOT A1 AND A0 AND B3 AND NOT B1 AND NOT B0) OR (A2 AND NOT A0
     AND NOT B2 AND B1 AND NOT B0) OR (NOT A2 AND A1 AND NOT A0 AND B2 AND NOT B0) OR (A3 AND NOT B3 AND NOT B2 AND NOT B1 AND B0) OR (NOT A3 AND A0 AND B3
     AND NOT B2 AND NOT B1) OR (A3 AND NOT A1 AND NOT A0 AND NOT B1 AND B0) OR (NOT A3 AND A2 AND NOT A1 AND A0 AND NOT B3 AND B2 AND NOT B1 AND B0) OR (
    NOT A3 AND NOT A2 AND A1 AND NOT B3 AND B2 AND NOT B1) OR (NOT A3 AND A2 AND NOT A1 AND NOT B3 AND NOT B2 AND B1) OR (NOT A3 AND NOT A2 AND A1 AND A0 AND NOT B3
     AND NOT B2 AND B1 AND B0) OR (A3 AND NOT A2 AND NOT A1 AND NOT A0 AND B0) OR (A2 AND NOT A1 AND NOT A0 AND B1 AND NOT B0) OR (A3 AND NOT A2 AND A1
     AND A0 AND B3 AND B2 AND NOT B1 AND B0) OR (NOT A3 AND A2 AND A1 AND A0 AND B3 AND B0) OR (A3 AND A2 AND NOT A1 AND A0 AND B3 AND NOT B2 AND B1 AND B0) OR (
    A3 AND A0 AND NOT B3 AND B2 AND B1 AND B0);

S2 <= (A2 AND A0 AND NOT B2 AND B0) OR (NOT A2 AND A0 AND B2 AND B0) OR (A0 AND B2 AND NOT B1 AND NOT B0) OR (A1 AND NOT B2 AND B1 AND NOT B0) OR (
    NOT A2 AND A1 AND NOT A0 AND B1) OR (A2 AND NOT A1 AND NOT A0 AND B0) OR (A1 AND NOT A0 AND B1 AND NOT B0) OR (NOT A1 AND A0 AND B2 AND NOT B0) OR (
    A2 AND NOT A0 AND NOT B1 AND B0);

S1 <= (A0 AND B1 AND NOT B0) OR (A1 AND NOT B1 AND B0) OR (A1 AND NOT A0 AND B0) OR (NOT A1 AND A0 AND B1);

S0 <= (A0 AND B0);

END data_flow;
