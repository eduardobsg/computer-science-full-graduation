LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY contador_primos IS
PORT (
	S5 : IN std_logic;
	S4 : IN std_logic;
	S3 : IN std_logic;
	S2 : IN std_logic;
	S1 : IN std_logic;
	S0 : IN std_logic;
	T5 : OUT std_logic;
	T4 : OUT std_logic;
	T3 : OUT std_logic;
	T2 : OUT std_logic;
	T1 : OUT std_logic;
	T0 : OUT std_logic);
END contador_primos;

ARCHITECTURE data_flow OF contador_primos IS
BEGIN

T5 <= (S5 AND S4 AND S3 AND S2 AND NOT S1 AND S0) OR(NOT S5 AND S4 AND S3 AND S2 AND S1 AND S0);

T4 <= (NOT S5 AND NOT S4 AND S3 AND S2 AND NOT S1 AND S0) OR(S5 AND S4 AND S3 AND S2 AND NOT S1 AND S0) OR(S5 AND NOT S4 AND S3 AND S2 AND S1 AND S0) OR(
    NOT S5 AND S4 AND S3 AND S2 AND S1 AND S0);

T3 <= (S5 AND NOT S3 AND S2 AND NOT S1 AND S0) OR(NOT S5 AND NOT S4 AND S3 AND S2 AND NOT S1 AND S0) OR(S5 AND S4 AND S2 AND NOT S1 AND S0) OR(
    NOT S5 AND NOT S3 AND S2 AND S1 AND S0) OR(S5 AND NOT S4 AND S3 AND S2 AND S1 AND S0) OR(NOT S5 AND S4 AND S2 AND S1 AND S0);

T2 <= (NOT S4 AND S3 AND NOT S2 AND S1 AND S0) OR(S5 AND S4 AND S2 AND NOT S1 AND S0) OR(S5 AND NOT S3 AND S2 AND NOT S1 AND S0) OR(NOT S5
     AND NOT S4 AND S3 AND S2 AND NOT S1 AND S0) OR(NOT S5 AND NOT S3 AND NOT S2 AND S1 AND S0) OR(S5 AND S3 AND NOT S2 AND S1 AND S0) OR(NOT S5
     AND NOT S4 AND NOT S3 AND S1 AND S0);

T1 <= (S4 AND S3 AND S2 AND NOT S1 AND S0) OR(NOT S5 AND NOT S4 AND NOT S3 AND NOT S2 AND NOT S1 AND NOT S0) OR(S5 AND NOT S4 AND S3 AND NOT S2 AND NOT S1
     AND S0) OR(S5 AND S4 AND S3 AND NOT S2 AND S1 AND S0) OR(S5 AND NOT S4 AND S3 AND S2 AND S1 AND S0) OR(S5 AND S4 AND S2 AND NOT S1 AND S0) OR(
    NOT S5 AND NOT S4 AND NOT S2 AND S1 AND S0) OR(NOT S5 AND S4 AND NOT S3 AND NOT S2 AND NOT S1 AND S0) OR(NOT S5 AND NOT S4 AND NOT S3 AND S2 AND NOT S1 AND S0) OR(
    NOT S5 AND S4 AND S2 AND S1 AND S0);

T0 <= (NOT S5 AND NOT S4 AND NOT S3 AND NOT S2 AND S1 AND NOT S0) OR(S5 AND S4 AND S3 AND S2 AND NOT S1 AND S0);

END data_flow;
